`include "d1.v"
`include "d2.v"
`include "dr.v"

module tia_audio_clock_divider(hphi1, hphi2, rhs, cnt, rcb, shs, lrhb, rsynl,
    rsynd, resphi0, hs, aphi1, aphi2
